
class MODULE_REGMAP;
endclass


